library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package typing_speed_pkg is
    constant CLOCK_FREQ : integer := 100_000; 
end package;